/****************************************************************************
 * axi4_2x2_uvm_env_pkg.sv
 ****************************************************************************/

/**
 * Package: axi4_2x2_uvm_env_pkg
 * 
 * TODO: Add package documentation
 */
`include "uvm_macros.svh" 
package axi4_2x2_uvm_env_pkg;
	import uvm_pkg::*;
	import axi4_master_agent_agent_pkg::*;
	
	`include "axi4_2x2_uvm_env.svh"

endpackage

