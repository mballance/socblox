
`include "uvm_macros.svh"

package axi4_uvm_master_agent_pkg;
	import uvm_pkg::*;
	
	`include "axi4_uvm_master_config.svh"
	`include "axi4_uvm_master_seq_item.svh"
	`include "axi4_uvm_master_driver.svh"
	`include "axi4_uvm_master_monitor.svh"
	`include "axi4_uvm_master_seq_base.svh"
	`include "axi4_uvm_master_agent.svh"
endpackage



